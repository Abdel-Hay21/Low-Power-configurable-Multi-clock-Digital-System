

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 8.373 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.2741 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 28.148 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 135.584 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.026 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.4175 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 221.322 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1070.82 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA45 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 5.225 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.1323 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 36.184 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 174.237 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 14.126 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.1385 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 283.123 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1368.09 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA45 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 1.981 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.52861 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 15.839 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.378 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.21 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 54.1125 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 220.984 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1069.2 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 1.456 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.19576 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 29.9372 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 146.956 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA23 ;
  END SI[0]
  PIN SO[3] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 3.626 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6335 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 47.4181 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 232.95 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 3.62207 LAYER VIA34 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 2.369 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.3949 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.00048 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.537 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.55 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 132.9 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 302.871 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1465 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.01839 LAYER VIA56 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 13.548 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1659 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.475 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.28715 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 23.629 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 113.848 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 158.989 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 768.131 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.30108 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 4.908 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.6075 LAYER METAL3 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.468 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.44348 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.65464 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.949327 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 4.71201 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 1.617 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77777 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.506 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 51.1111 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 96.8762 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 475.143 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.37054 LAYER VIA45 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 2.993 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3963 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 14.922 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.1596 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6822 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 39.9929 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 194.032 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.076 LAYER VIA45 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 2.041 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.81721 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.361 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3588 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.1145 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 122.218 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA34 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 6.235 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1828 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.937 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3194 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 60.8443 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 296.415 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.3546 LAYER VIA34 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.269 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29389 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.41558 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.00287 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 4.96957 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.301 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.44781 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.258 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.9134 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.733512 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 3.67394 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 7.639 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.7436 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 19.952 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.3539 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6162 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 50.6502 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 243.475 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.527264 LAYER VIA34 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNAPARTIALMETALAREA 5.053 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.3049 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNADIFFAREA 1.529 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 6.573 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.8085 LAYER METAL4 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 2.515 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0972 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 20.531 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 98.9465 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3328 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 91.6003 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 445.88 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.70016 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 2.447 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7701 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 22.08 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 106.397 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4108 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 69.6063 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 336.141 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.878773 LAYER VIA56 ;
  END framing_error
END SYS_TOP

END LIBRARY
